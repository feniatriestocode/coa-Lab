`include "constants.h"

/************** Main control in ID pipe stage  *************/
module control_main(output reg RegDst,
                output reg Branch,  
                output reg MemRead,
                output reg MemWrite,  
                output reg MemToReg,  
                output reg ALUSrc,  
                output reg RegWrite,  
                output reg BneEn,  
                output reg [1:0] ALUcntrl,  
                input [5:0] opcode);

  always @(*) 
   begin
     case (opcode)
      `R_FORMAT: 
      /* TO FILL IN: The control signal values in each and every case */
          begin 
            RegDst 		= 1'b1;
            MemRead 	= 1'b0;
            MemWrite 	= 1'b0;
            MemToReg 	= 1'b0;
            ALUSrc 		= 1'b0;
            Branch 		= 1'b0;     
            ALUcntrl 	= 2'b10;
			BneEn		= 1'b1;
            #(`clock_period / 4) RegWrite = 1'b1;
            #(`clock_period / 2) RegWrite = 1'b0;
          end
       `LW :   
           begin 
            RegDst 		= 1'b1;
            MemRead 	= 1'b0;
            MemWrite 	= 1'b0;
            MemToReg 	= 1'b0;
            ALUSrc 		= 1'b0;
            Branch 		= 1'b0;     
            ALUcntrl 	= 2'b10;            
            #(`clock_period / 4) RegWrite = 1'b1;
            #(`clock_period / 2) RegWrite = 1'b0;
           end
        `SW :   
           begin 
            RegDst 		= 1'b1;
            MemRead 	= 1'b0;
            MemWrite 	= 1'b0;
            MemToReg 	= 1'b0;
            ALUSrc 		= 1'b0;
            Branch 		= 1'b0;     
            ALUcntrl 	= 2'b10;            
            #(`clock_period / 4) RegWrite = 1'b1;
            #(`clock_period / 2) RegWrite = 1'b0;
           end
       `BEQ:  
           begin 
            RegDst 		= 1'b1;
            MemRead 	= 1'b0;
            MemWrite 	= 1'b0;
            MemToReg 	= 1'b0;
            ALUSrc 		= 1'b0;
            Branch 		= 1'b0;     
            ALUcntrl 	= 2'b10;            
            #(`clock_period / 4) RegWrite = 1'b1;
            #(`clock_period / 2) RegWrite = 1'b0;
           end
       default:
           begin
            RegDst 		= 1'b0;
            MemRead 	= 1'b0;
            MemWrite 	= 1'b0;
            MemToReg 	= 1'b0;
            ALUSrc 		= 1'b0;
            Branch 		= 1'b0;     
            ALUcntrl 	= 2'b00;            
            RegWrite = 1'b0;
           end
      endcase
    end // always
endmodule


/**************** Module for Bypass Detection in EX pipe stage goes here  *********/
// TO FILL IN: Module details 
endmodule          
                       

/**************** Module for Stall Detection in ID pipe stage goes here  *********/
// TO FILL IN: Module details 

                       
/************** control for ALU control in EX pipe stage  *************/
module control_alu(output reg [3:0] ALUOp,                  
               input [1:0] ALUcntrl,
               input [5:0] func);

  always @(ALUcntrl or func)  
    begin
      case (ALUcntrl)
        2'b10: 
           begin
             case (func)
              6'b100000: ALUOp  = 4'b0010; // add
              6'b100010: ALUOp = 4'b0110; // sub
              6'b100100: ALUOp = 4'b0000; // and
              6'b100101: ALUOp = 4'b0001; // or
              6'b100111: ALUOp = 4'b1100; // nor
              6'b101010: ALUOp = 4'b0111; // slt
              default: ALUOp = 4'b0000;       
             endcase 
          end   
        2'b00: 
              ALUOp  = 4'b0010; // add
        2'b01: 
              ALUOp = 4'b0110; // sub
        default:
              ALUOp = 4'b0000;
     endcase
    end
endmodule
